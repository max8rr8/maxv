

`default_nettype none

module code (
    input clk_i,
    input [31:0] addr_i,
    output [31:0] instr_o
);
  pROM #(
    .BIT_WIDTH(16),
.INIT_RAM_00(256'b0000000000000000000000000110111100000000010101010000000000100011000001101001000000000010100100111111111000000011000111101110001111111111111100110000001100010011000000000000000000100011001101110000000001010101000000000010001100000110000100000000001010010011),
.INIT_RAM_01(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000110111100000000000000000000000001101111),
.INIT_RAM_02(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_03(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_04(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_05(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_06(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_07(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_08(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_09(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_0A(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_0B(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_0C(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_0D(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_0E(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_0F(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_10(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_11(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_12(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_13(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_14(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_15(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_16(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_17(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_18(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_19(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_1A(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_1B(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_1C(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_1D(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_1E(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_1F(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_20(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_21(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_22(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_23(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_24(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_25(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_26(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_27(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_28(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_29(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_2A(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_2B(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_2C(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_2D(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_2E(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_2F(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_30(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_31(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_32(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_33(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_34(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_35(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_36(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_37(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_38(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_39(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_3A(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_3B(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_3C(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_3D(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_3E(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_3F(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),

    .READ_MODE(0),
    .RESET_MODE("SYNC")
  ) prom_inst_lo (
      .AD({addr_i[11:0], 2'b0}),
      .CE(1'b1),
      .CLK(clk_i),
      .DO(instr_o[15:0]),
      .OCE(1'b1),
      .RESET(1'b0)
  );

	pROM #(
    .BIT_WIDTH(16),
.INIT_RAM_00(256'b0000000000000000000000000110111100000000010101010000000000100011000001101001000000000010100100111111111000000011000111101110001111111111111100110000001100010011000000000000000000100011001101110000000001010101000000000010001100000110000100000000001010010011),
.INIT_RAM_01(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000110111100000000000000000000000001101111),
.INIT_RAM_02(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_03(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_04(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_05(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_06(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_07(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_08(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_09(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_0A(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_0B(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_0C(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_0D(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_0E(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_0F(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_10(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_11(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_12(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_13(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_14(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_15(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_16(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_17(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_18(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_19(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_1A(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_1B(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_1C(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_1D(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_1E(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_1F(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_20(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_21(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_22(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_23(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_24(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_25(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_26(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_27(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_28(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_29(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_2A(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_2B(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_2C(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_2D(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_2E(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_2F(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_30(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_31(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_32(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_33(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_34(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_35(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_36(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_37(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_38(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_39(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_3A(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_3B(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_3C(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_3D(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_3E(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),
.INIT_RAM_3F(256'b0000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011000000000000000000000000000100110000000000000000000000000001001100000000000000000000000000010011),

    .READ_MODE(0),
    .RESET_MODE("SYNC")
  ) prom_inst_hi (
      .AD({addr_i[11:0], 2'b0}),
      .CE(1'b1),
      .CLK(clk_i),
      .DO(instr_o[31:16]),
      .OCE(1'b1),
      .RESET(1'b0)
  );
endmodule
