
  package vde_init_mem;
    localparam logic [55299:0] MEM_MAP_INIT = 'h7fbfc00ff00001fe00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003fdfe007f801fe000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007f801fe00003fdfe00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004048a0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000404880000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000404ac00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    localparam logic [65535:0] MEM_SPRITE_INIT = 65536'h6040200000000008000000080003c008000787080006c788000ec0f8000180080001800800000388000760080000030800018188000180e800018188000606080003030800000008000cc788000c0388000db068000db008000cc1c80006c388000c6388000ccfc80001800800066008000d800800060fc80006c008000c0008000cc008000c800800000ff80000f0f8000f0f08000ff008000ffff80001f008000f8188000ff188000ff3680003f0080001f0080001f1880003f368000ff008000ff008000ff368000ff188000f7368000ff00800037368000f7008000ff368000370080003f368000373680001f188000ff188000ff0080001f188000ff008000ff1880001f188000f8008000f8188000fe368000fe368000f600800036368000f6368000f8008000fe008000f6368000f8188000f818800018188000dbdb8000555580002222800066008000660080001818800037c3800033c380000c008000c0008000c030800000388000003c8000fcfc8000cc008000cc008000cc008000303880007c1c8000180e8000c6f8800030cc800060388000c0188000cccc800066c38000cc008000cc008000cc788000cc008000cc008000cc788000cc3e80007f008000781c8000cc308000fec6800030e08000187c800030cc8000fce08000fccc80007e7e8000c00080007c3080007ce080007ccc80003e7e8000fc1c8000cc00800078788000c60080000076800030e0800018188000301c800030008000cc00800038008000fe008000cc008000cc008000301080007800800066008000cc00800066008000cc008000cc008000fe0080003070800078e080000c0c80003030800066e08000cc00800060388000fc008000cc1c8000c000800066e080007c008000003080000000800000108000187880000cc080006078800032fe800030cc800038c68000fec68000cccc8000cccc800030fc80001c7880006cfc8000dc78800060fc8000c6388000cec68000d6c6800062f080006ce68000cc1e800030788000cccc8000ce3c800068fe800068fe800066f88000c03c800066fc8000fc308000de7c80003078800018608000000080006018800000008000000080000c788000cc78800030fc8000cc3880000cfc8000fe1c80000c7880006078800030308000f67c800060068000000080000000800000008000300080003c008000186080006018800000608000dc388000300080000c308000fe6c8000006c800030308000000080003c008000ff00800066008000c0008000600080000c0080007e188000181880007e1880007e0080006c3e80001b7f800066668000181880003e028000f8808000e7998000637f8000303f80003c3c8000cc0f8000bdff800042008000c3ff80003c008000fe108000fe3880007c1080007c6c8000c37e8000bd7e80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007050301000000000000000000003c00000000180000006c00006c0c00000000000000000000006c0000dc76000030300000d8180000181b0000003000000030000000300000fcfc0000cccc0000606000007e0c00007e000000cc3000006c6c00006c6c000078300000187600007c660000d8000000cccc00006cfe0000c0fc0000f8780000dc00000000ff00000f0f0000f0f00000ff000000ffff00001800000000180000181800003636000036000000180000000018000000360000360000001800000000360000001800003636000000000000363600003600000000360000360000000036000036360000181800001818000000000000181800001800000000180000001800001800000000180000003600000036000036000000363600003636000018000000360000003636000018180000181800001818000077770000aaaa000088880000cccc000033330000181800006fc6000066c600000c000000c0000000cc0000007c6c00007e6c0000dc000000ccf80000cc1c0000cc1c000030000000cc000000181b0000cfcc0000fccc0000e66c00007e180000cc0000003c1800007ccc0000cce00000cccc0000cce00000cccc0000cccc0000cc6c0000cc00000060000000fc300000c63800003000000018c6000030000000c0000000c000000060c3000078000000cc300000cc000000cc00000066c30000c0000000cccc000018cc0000c610000000dc0000303000001818000030300000640000007c0000006c000000fe00000078000000cc000000343000000c000000600000007c0000007c000000cc000000cc000000d6000000303000006c600000cc00000030000000666000007c000000606c0000c0000000cc0c0000cc00000066600000cc00000000300000000000000038000018180000066000006060000066c6000030cc00006cc60000eec6000078cc0000cccc000030b40000cccc00006666000078cc0000606600006c6c0000c6e60000c6ee00006660000066660000cc0c000030300000cccc00006666000060620000626200006c6c00006666000066660000cc780000c0c6000000cc000030300000fc00000030300000303000003030000018cc0000cccc000030cc0000cc600000ccc000000c3c0000cccc0000cccc000030700000e6c60000c00c00003000000000000000300000003030000066660000303000003030000000600000cc6c000066c60000f87c00006c6c0000006c0000007800000000000018ff0000ff18000024240000fe00000030300000181800003c180000183c00003c3c00007e000000386300001bdb0000006600007e3c00000e0e0000e0e000003c5a0000676300007033000018660000cc07000099c30000663c0000e7ff0000180000007c1000007c7c00003838000038fe0000e7ff000099810000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006040200000000010000000100003c010000300100006c01003c0c01000000010000000100006c010000dc010030000100d8180100181b0100fc600100fc180100fcfc010000000100cccc010038c00100607e0100007e010078180100eec6010038c601003078010018dc010060660100707e0100fc6001006c6c0100c0cc0100c0cc01007676010000ff01000f0f0100f0f00100ff000100ffff0100180001000018010018ff01003636010036000100181f0100001f0100003601003600010018ff01000036010000ff010036f7010000ff01003637010036ff010000f70100363f01000037010036360100181f01001818010000000100181801001800010000180100001801001800010000f801000036010000f6010036fe01003636010036f6010018f80100360001003636010018f801001818010018180100dbdb01005555010022220100006601000066010018000100cfcc0100cccc0100000001000000010078300100006c0100006c0100cccc0100cc0001007e00010078000100787001007e780100d8180100c6cc010030780100fc640100187e010078cc0100183c01000c0001007e0001007e000100780001007800010078000100cecc01007f7f0100fcfc0100cc000100c66c0100787001003c3801007870010078780100787801003c3c01000c7801007e7801007e7801007e7801003f3c0100787801007e0001000cc00100fe38010000000100e0300100181801001c300100fcfc01000ccc0100c6c601006cc6010030cc010076cc0100187c0100f87c0100f0dc01000c76010060dc010078780100ccf80100c6cc010078300100e6660100cc0c010078700100e66c01000c760100f060010078780100760c010078780100dc600100767801000018010000000100006c0100781801000230010078600100fe8c010078cc0100c66c0100c6c6010030cc0100fccc01007830010078e00100e66601001ccc0100f066010038c60100c6f60100c6fe0100fe600100e66c0100780c010078300100cccc01003ec00100f0680100fe680100f86601003cc00100fc660100cccc010078de0100300c01006018010000fc010018600100303001003030010070cc010078cc0100300c010078c0010078f801001e6c0100780c0100fc0c0100fc3001007cce01008018010030000100000001003000010000300100003c0100601801001860010000c0010076380100c6cc010030c001006cfe0100006c0100307801000000010000ff0100003c01000066010000c0010000600100000c010018180100187e0100187e01007e000100cc3801001bdb0100666601003c7e0100023e010080f801005a3c0100e67f0100f03f01007e660100cc0f0100c39901003c660100ffe70100001801003838010038380100107c010010fe0100ffdb010081a50100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000107050300000000000000000000003c000000600000006c00001c0c00000000000000180000003800000000000000fc0000701800001818000000300000003000000030000000fc000000cc000000f80000c0db000000db0000007c000000c6000000fe0000fccc000000180000c066000000d8000000300000006c000000c00000c0f8000000dc000000ff00000f0f0000f0f00000ff000000ffff000018000000001800001818000036360000360000001818000000180000003600003600000018000000003600000000000036000000000000003630000036000000000000003630000000300000363600001818000018180000000000001818000018000000001800000018000018000000001800000036000000060000360600003636000036060000181800003600000036360000181800001818000018180000eeee0000aaaa0000888800000033000000cc00000018000003db00000fde000000fc000000fc00000060000000380000003e000000ec000000f8000000cc00000078000000300000000c0000703c0000c7fa000030fc000000f0000018c0000000cc000000660000f8cc000000cc000000cc000000780000007800000078000000fe0000000c0000006000000078000000c6000000300000001800000030000000cc000000cc00000066000038c00000000c0000000c0000000c00000006000000cc000000cc000078cc0000006c000000000000001c00000000000000e0000000980000f8cc0000006c000000d6000000cc000000cc00000030000000c00000007600001ecc0000f066000000cc000000cc000000fe000000300000006c0000780c00000030000000760000f8cc000000f0000000cc0000007c000000cc0000007c0000000c000000000000ff00000000c6000000180000001800000060000000180000007800000038000000d6000000cc000000cc00000030000000700000007c000000cc0000007c000000c6000000de000000fe00000060000000780000000c00000030000000fc000000c0000000780000007800000066000000c00000007c000000cc000000de000000180000000c00000000000000c000006000000000000000007c0000007800000018000000f80000000c000000cc000000380000003800000030000000de0000003000000000000000fc00006000000000fc000000ff0000001800000060000000000000007600000018000000780000006c0000000000000030000000000000007e0000007e000000ff000000c0000000fe000000fe00000018000000180000ff18000000000000786c0000007b0000006600001818000000fe000000fe000099e70000c0630000e030000018660000787d0000ffbd000000420000ffc30000003c00007c7c00007cfe000000fe000000fe00007eff00007e8100000000;
  endpackage
  