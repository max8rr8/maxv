//Credit to the Implementation of HDMI Spec v1.4a by Sameer Puri https://github.com/sameer
`default_nettype none

module dvi_pattern (
    input wire clk_i,
    input logic rstn_i,

    // Pixel input
    input wire [23:0] display_data_i,
    input wire display_valid_i,
    output wire display_ready_o,
    output wire display_clk_o,

    // Frame track
    output wire frame_toggle_o,

    // HDMI Output
    output wire tmds_clk_n_o,
    output wire tmds_clk_p_o,
    output wire [2:0] tmds_d_n_o,
    output wire [2:0] tmds_d_p_o,
);
  wire clk_pixel, clk_display_x5, pll_lock, reset;
  logic [2:0] tmds;
  logic       tmds_clock;

  assign reset = ~rstn_i;

  PLL480 pll_dvi (
      .clkin (clk_i),
      .clkout(clk_display_x5),
      .lock  (pll_lock)
  );

  CLKDIV #(
      .DIV_MODE("5")
  ) clk_div (
      .CLKOUT(clk_pixel),
      .HCLKIN(clk_display_x5),
      .RESETN(pll_lock)
  );

  assign display_clk_o = clk_pixel;


  localparam BIT_WIDTH = 10;
  localparam BIT_HEIGHT = 10;
  localparam START_X = 0;
  localparam START_Y = 0;
  localparam int NUM_CHANNELS = 3;
  logic hsync;
  logic vsync;

  logic [BIT_WIDTH-1:0] cx = START_X;
  logic [BIT_HEIGHT-1:0] cy = START_Y;


  localparam real VIDEO_RATE = 25.2E6;

  localparam [BIT_WIDTH-1:0] FRAME_WIDTH = 800;
  localparam [BIT_HEIGHT-1:0] FRAME_HEIGHT = 525;
  localparam [BIT_WIDTH-1:0] SCREEN_WIDTH = 640;
  localparam [BIT_HEIGHT-1:0] SCREEN_HEIGHT = 480;
  localparam [BIT_WIDTH-1:0] HSYNC_PULSE_START = 16;
  localparam [BIT_WIDTH-1:0] HSYNC_PULSE_SIZE = 96;
  localparam [BIT_HEIGHT-1:0] VSYNC_PULSE_START = 10;
  localparam [BIT_HEIGHT-1:0] VSYNC_PULSE_SIZE = 2;
  localparam INVERT = 1;


  wire next = screen_partition == (SCREEN_WIDTH - 1'B1);
  reg [BIT_WIDTH-1:0] screen_partition;

  reg [23:0] old_color, new_color;

  always_comb begin
    hsync <= INVERT ^ (cx >= SCREEN_WIDTH + HSYNC_PULSE_START && cx < SCREEN_WIDTH + HSYNC_PULSE_START + HSYNC_PULSE_SIZE);
    // vsync pulses should begin and end at the start of hsync, so special
    // handling is required for the lines on which vsync starts and ends
    if (cy == SCREEN_HEIGHT + VSYNC_PULSE_START)
      vsync <= INVERT ^ (cx >= SCREEN_WIDTH + HSYNC_PULSE_START);
    else if (cy == SCREEN_HEIGHT + VSYNC_PULSE_START + VSYNC_PULSE_SIZE)
      vsync <= INVERT ^ (cx < SCREEN_WIDTH + HSYNC_PULSE_START);
    else
      vsync <= INVERT ^ (cy >= SCREEN_HEIGHT + VSYNC_PULSE_START && cy < SCREEN_HEIGHT + VSYNC_PULSE_START + VSYNC_PULSE_SIZE);
  end

  // Wrap-around pixel position counters indicating the pixel to be generated by the user in THIS clock and sent out in the NEXT clock.
  always_ff @(posedge clk_pixel) begin
    if (reset) begin
      cx <= BIT_WIDTH'(START_X);
      cy <= BIT_HEIGHT'(START_Y);
    end else begin
      cx <= cx == FRAME_WIDTH - 1'b1 ? BIT_WIDTH'(0) : cx + 1'b1;
      cy <= cx == FRAME_WIDTH - 1'b1 ? cy == FRAME_HEIGHT - 1'b1 ? BIT_HEIGHT'(0) : cy + 1'b1 : cy;
    end
  end

  always_ff @(posedge clk_pixel) begin
    if(reset) begin
        frame_toggle_o <= 0;
    end else begin
        if(cy == SCREEN_HEIGHT && cx == 0) begin
            frame_toggle_o <= ~frame_toggle_o;
        end
    end
  end

  // See Section 5.2
  logic video_data_period = 0;
  always_ff @(posedge clk_pixel) begin
    if (reset) video_data_period <= 0;
    else video_data_period <= cx < SCREEN_WIDTH && cy < SCREEN_HEIGHT;
  end

  assign display_ready_o = video_data_period;

  logic [ 2:0] mode = 3'd1;
  logic [23:0] video_data = 24'd0;
  logic [ 5:0] control_data = 6'd0;
  logic [11:0] data_island_data = 12'd0;

  always_ff @(posedge clk_pixel) begin
    if (reset) begin
      mode <= 3'd0;
      video_data <= 24'd0;
      control_data <= 6'd0;
    end else begin
      mode <= video_data_period ? 3'd1 : 3'd0;
      video_data <= display_data_i;
      control_data <= {4'b0000, {vsync, hsync}};  // ctrl3, ctrl2, ctrl1, ctrl0, vsync, hsync
    end
  end


  // All logic below relates to the production and output of the 10-bit TMDS code.
  logic [9:0] tmds_internal[NUM_CHANNELS-1:0]  /* verilator public_flat */;
  genvar i;
  generate
    // TMDS code production.
    for (i = 0; i < NUM_CHANNELS; i++) begin : tmds_gen
      tmds_channel #(
          .CN(i)
      ) tmds_channel (
          .clk_pixel(clk_pixel),
          .video_data(video_data[i*8+7:i*8]),
          .data_island_data(0),
          .control_data(control_data[i*2+1:i*2]),
          .mode(mode),
          .tmds(tmds_internal[i])
      );
    end
  endgenerate


  OSER10 gwSer0 (
      .Q(tmds[0]),
      .D0(tmds_internal[0][0]),
      .D1(tmds_internal[0][1]),
      .D2(tmds_internal[0][2]),
      .D3(tmds_internal[0][3]),
      .D4(tmds_internal[0][4]),
      .D5(tmds_internal[0][5]),
      .D6(tmds_internal[0][6]),
      .D7(tmds_internal[0][7]),
      .D8(tmds_internal[0][8]),
      .D9(tmds_internal[0][9]),
      .PCLK(clk_pixel),
      .FCLK(clk_display_x5),
      .RESET(reset)
  );

  OSER10 gwSer1 (
      .Q(tmds[1]),
      .D0(tmds_internal[1][0]),
      .D1(tmds_internal[1][1]),
      .D2(tmds_internal[1][2]),
      .D3(tmds_internal[1][3]),
      .D4(tmds_internal[1][4]),
      .D5(tmds_internal[1][5]),
      .D6(tmds_internal[1][6]),
      .D7(tmds_internal[1][7]),
      .D8(tmds_internal[1][8]),
      .D9(tmds_internal[1][9]),
      .PCLK(clk_pixel),
      .FCLK(clk_display_x5),
      .RESET(reset)
  );

  OSER10 gwSer2 (
      .Q(tmds[2]),
      .D0(tmds_internal[2][0]),
      .D1(tmds_internal[2][1]),
      .D2(tmds_internal[2][2]),
      .D3(tmds_internal[2][3]),
      .D4(tmds_internal[2][4]),
      .D5(tmds_internal[2][5]),
      .D6(tmds_internal[2][6]),
      .D7(tmds_internal[2][7]),
      .D8(tmds_internal[2][8]),
      .D9(tmds_internal[2][9]),
      .PCLK(clk_pixel),
      .FCLK(clk_display_x5),
      .RESET(reset)
  );

  assign tmds_clock = clk_pixel;

  ELVDS_OBUF tmds_bufds[3:0] (
      .I ({clk_pixel, tmds}),
      .O ({tmds_clk_p_o, tmds_d_p_o}),
      .OB({tmds_clk_n_o, tmds_d_n_o})
  );
endmodule
